
module Nios2Computer (
	clk_clk,
	led_pio_ext_connection_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	led_pio_ext_connection_export;
	input		reset_reset_n;
endmodule
